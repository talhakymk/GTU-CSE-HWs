module mux_and(output [31:0] res ,input [31:0] a, input [31:0] b , input [31:0] c , input [31:0] d);
	and(res[0] , a[0] , b[0] , c[0] , d[0]);
	and(res[1] , a[1] , b[1] , c[1] , d[1]);
	and(res[2] , a[2] , b[2] , c[2] , d[2]);
	and(res[3] , a[3] , b[3] , c[3] , d[3]);
	and(res[4] , a[4] , b[4] , c[4] , d[4]);
	and(res[5] , a[5] , b[5] , c[5] , d[5]);
	and(res[6] , a[6] , b[6] , c[6] , d[6]);
	and(res[7] , a[7] , b[7] , c[7] , d[7]);
	and(res[8] , a[8] , b[8] , c[8] , d[8]);
	and(res[9] , a[9] , b[9] , c[9] , d[9]);
	and(res[10] , a[10] , b[10] , c[10] , d[10]);
	and(res[11] , a[11] , b[11] , c[11] , d[11]);
	and(res[12] , a[12] , b[12] , c[12] , d[12]);
	and(res[13] , a[13] , b[13] , c[13] , d[13]);
	and(res[14] , a[14] , b[14] , c[14] , d[14]);
	and(res[15] , a[15] , b[15] , c[15] , d[15]);
	and(res[16] , a[16] , b[16] , c[16] , d[16]);
	and(res[17] , a[17] , b[17] , c[17] , d[17]);
	and(res[18] , a[18] , b[18] , c[18] , d[18]);
	and(res[19] , a[19] , b[19] , c[19] , d[19]);
	and(res[20] , a[20] , b[20] , c[20] , d[20]);
	and(res[21] , a[21] , b[21] , c[21] , d[21]);
	and(res[22] , a[22] , b[22] , c[22] , d[22]);
	and(res[23] , a[23] , b[23] , c[23] , d[23]);
	and(res[24] , a[24] , b[24] , c[24] , d[24]);
	and(res[25] , a[25] , b[25] , c[25] , d[25]);
	and(res[26] , a[26] , b[26] , c[26] , d[26]);
	and(res[27] , a[27] , b[27] , c[27] , d[27]);
	and(res[28] , a[28] , b[28] , c[28] , d[28]);
	and(res[29] , a[29] , b[29] , c[29] , d[29]);
	and(res[30] , a[30] , b[30] , c[30] , d[30]);
	and(res[31] , a[31] , b[31] , c[31] , d[31]);
endmodule
	