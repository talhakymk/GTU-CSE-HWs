module full_adder(output r,p,g , input a , b , c_in);
	
endmodule
